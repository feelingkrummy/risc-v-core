module decode (

);

endmodule
